magic
tech gf180mcuD
magscale 1 10
timestamp 1702315505
<< nwell >>
rect 1258 235552 558742 236416
rect 1258 233984 558742 234848
rect 1258 232416 558742 233280
rect 1258 230848 558742 231712
rect 1258 229280 558742 230144
rect 1258 227712 558742 228576
rect 1258 226144 558742 227008
rect 1258 224576 558742 225440
rect 1258 223008 558742 223872
rect 1258 221440 558742 222304
rect 1258 219872 558742 220736
rect 1258 218304 558742 219168
rect 1258 216736 558742 217600
rect 1258 215168 558742 216032
rect 1258 213600 558742 214464
rect 1258 212032 558742 212896
rect 1258 210464 558742 211328
rect 1258 208896 558742 209760
rect 1258 207328 558742 208192
rect 1258 205760 558742 206624
rect 1258 204192 558742 205056
rect 1258 202624 558742 203488
rect 1258 201056 558742 201920
rect 1258 199488 558742 200352
rect 1258 197920 558742 198784
rect 1258 196352 558742 197216
rect 1258 194784 558742 195648
rect 1258 193216 558742 194080
rect 1258 191648 558742 192512
rect 1258 190080 558742 190944
rect 1258 188512 558742 189376
rect 1258 186944 558742 187808
rect 1258 185376 558742 186240
rect 1258 183808 558742 184672
rect 1258 182240 558742 183104
rect 1258 180672 558742 181536
rect 1258 179104 558742 179968
rect 1258 177536 558742 178400
rect 1258 175968 558742 176832
rect 1258 174400 558742 175264
rect 1258 172832 558742 173696
rect 1258 171264 558742 172128
rect 1258 169696 558742 170560
rect 1258 168128 558742 168992
rect 1258 166560 558742 167424
rect 1258 164992 558742 165856
rect 1258 163424 558742 164288
rect 1258 161856 558742 162720
rect 1258 160288 558742 161152
rect 1258 158720 558742 159584
rect 1258 157152 558742 158016
rect 1258 155584 558742 156448
rect 1258 154016 558742 154880
rect 1258 152448 558742 153312
rect 1258 150880 558742 151744
rect 1258 149312 558742 150176
rect 1258 147744 558742 148608
rect 1258 146176 558742 147040
rect 1258 144608 558742 145472
rect 1258 143040 558742 143904
rect 1258 141472 558742 142336
rect 1258 139904 558742 140768
rect 1258 138363 558742 139200
rect 1258 138336 276656 138363
rect 1258 137605 271392 137632
rect 1258 136795 558742 137605
rect 1258 136768 274752 136795
rect 1258 136039 273824 136064
rect 1258 136037 286176 136039
rect 1258 135227 558742 136037
rect 1258 135200 268144 135227
rect 1258 134471 287198 134496
rect 1258 134469 293568 134471
rect 1258 133632 558742 134469
rect 1258 132901 294128 132928
rect 1258 132091 558742 132901
rect 1258 132064 267696 132091
rect 1258 131333 265904 131360
rect 1258 130523 558742 131333
rect 1258 130496 281920 130523
rect 1258 129765 264336 129792
rect 1258 128955 558742 129765
rect 1258 128928 266128 128955
rect 1258 128197 286512 128224
rect 1258 127360 558742 128197
rect 1258 126629 265120 126656
rect 1258 125792 558742 126629
rect 1258 125061 264448 125088
rect 1258 124251 558742 125061
rect 1258 124224 285616 124251
rect 1258 122683 558742 123520
rect 1258 122656 266128 122683
rect 1258 121927 271805 121952
rect 1258 121925 301408 121927
rect 1258 121115 558742 121925
rect 1258 121088 267248 121115
rect 1258 119547 558742 120384
rect 1258 119520 301296 119547
rect 1258 118791 290402 118816
rect 1258 117977 558742 118791
rect 1258 117952 288766 117977
rect 1258 117221 273856 117248
rect 1258 116411 558742 117221
rect 1258 116384 275536 116411
rect 1258 115653 278336 115680
rect 1258 114843 558742 115653
rect 1258 114816 283040 114843
rect 1258 114085 271616 114112
rect 1258 113275 558742 114085
rect 1258 113248 268144 113275
rect 1258 112517 264448 112544
rect 1258 111680 558742 112517
rect 1258 110951 274542 110976
rect 1258 110949 277888 110951
rect 1258 110139 558742 110949
rect 1258 110112 284048 110139
rect 1258 109381 263664 109408
rect 1258 108571 558742 109381
rect 1258 108544 292560 108571
rect 1258 107815 276894 107840
rect 1258 107813 279344 107815
rect 1258 107003 558742 107813
rect 1258 106976 284608 107003
rect 1258 106245 264784 106272
rect 1258 105408 558742 106245
rect 1258 104677 270048 104704
rect 1258 103840 558742 104677
rect 1258 103109 277888 103136
rect 1258 102297 558742 103109
rect 1258 102272 278518 102297
rect 1258 100704 558742 101568
rect 1258 99136 558742 100000
rect 1258 97568 558742 98432
rect 1258 96000 558742 96864
rect 1258 94432 558742 95296
rect 1258 92864 558742 93728
rect 1258 91296 558742 92160
rect 1258 89728 558742 90592
rect 1258 88160 558742 89024
rect 1258 86592 558742 87456
rect 1258 85024 558742 85888
rect 1258 83456 558742 84320
rect 1258 81888 558742 82752
rect 1258 80320 558742 81184
rect 1258 78752 558742 79616
rect 1258 77184 558742 78048
rect 1258 75616 558742 76480
rect 1258 74048 558742 74912
rect 1258 72480 558742 73344
rect 1258 70912 558742 71776
rect 1258 69344 558742 70208
rect 1258 67776 558742 68640
rect 1258 66208 558742 67072
rect 1258 64640 558742 65504
rect 1258 63072 558742 63936
rect 1258 61504 558742 62368
rect 1258 59936 558742 60800
rect 1258 58368 558742 59232
rect 1258 56800 558742 57664
rect 1258 55232 558742 56096
rect 1258 53664 558742 54528
rect 1258 52096 558742 52960
rect 1258 50528 558742 51392
rect 1258 48960 558742 49824
rect 1258 47392 558742 48256
rect 1258 45824 558742 46688
rect 1258 44256 558742 45120
rect 1258 42688 558742 43552
rect 1258 41120 558742 41984
rect 1258 39552 558742 40416
rect 1258 37984 558742 38848
rect 1258 36416 558742 37280
rect 1258 34848 558742 35712
rect 1258 33280 558742 34144
rect 1258 31712 558742 32576
rect 1258 30144 558742 31008
rect 1258 28576 558742 29440
rect 1258 27008 558742 27872
rect 1258 25440 558742 26304
rect 1258 23872 558742 24736
rect 1258 22304 558742 23168
rect 1258 20736 558742 21600
rect 1258 19168 558742 20032
rect 1258 17600 558742 18464
rect 1258 16032 558742 16896
rect 1258 14464 558742 15328
rect 1258 12896 558742 13760
rect 1258 11328 558742 12192
rect 1258 9760 558742 10624
rect 1258 8192 558742 9056
rect 1258 6624 558742 7488
rect 1258 5056 558742 5920
rect 1258 3488 558742 4352
<< pwell >>
rect 1258 236416 558742 236854
rect 1258 234848 558742 235552
rect 1258 233280 558742 233984
rect 1258 231712 558742 232416
rect 1258 230144 558742 230848
rect 1258 228576 558742 229280
rect 1258 227008 558742 227712
rect 1258 225440 558742 226144
rect 1258 223872 558742 224576
rect 1258 222304 558742 223008
rect 1258 220736 558742 221440
rect 1258 219168 558742 219872
rect 1258 217600 558742 218304
rect 1258 216032 558742 216736
rect 1258 214464 558742 215168
rect 1258 212896 558742 213600
rect 1258 211328 558742 212032
rect 1258 209760 558742 210464
rect 1258 208192 558742 208896
rect 1258 206624 558742 207328
rect 1258 205056 558742 205760
rect 1258 203488 558742 204192
rect 1258 201920 558742 202624
rect 1258 200352 558742 201056
rect 1258 198784 558742 199488
rect 1258 197216 558742 197920
rect 1258 195648 558742 196352
rect 1258 194080 558742 194784
rect 1258 192512 558742 193216
rect 1258 190944 558742 191648
rect 1258 189376 558742 190080
rect 1258 187808 558742 188512
rect 1258 186240 558742 186944
rect 1258 184672 558742 185376
rect 1258 183104 558742 183808
rect 1258 181536 558742 182240
rect 1258 179968 558742 180672
rect 1258 178400 558742 179104
rect 1258 176832 558742 177536
rect 1258 175264 558742 175968
rect 1258 173696 558742 174400
rect 1258 172128 558742 172832
rect 1258 170560 558742 171264
rect 1258 168992 558742 169696
rect 1258 167424 558742 168128
rect 1258 165856 558742 166560
rect 1258 164288 558742 164992
rect 1258 162720 558742 163424
rect 1258 161152 558742 161856
rect 1258 159584 558742 160288
rect 1258 158016 558742 158720
rect 1258 156448 558742 157152
rect 1258 154880 558742 155584
rect 1258 153312 558742 154016
rect 1258 151744 558742 152448
rect 1258 150176 558742 150880
rect 1258 148608 558742 149312
rect 1258 147040 558742 147744
rect 1258 145472 558742 146176
rect 1258 143904 558742 144608
rect 1258 142336 558742 143040
rect 1258 140768 558742 141472
rect 1258 139200 558742 139904
rect 1258 137632 558742 138336
rect 1258 136064 558742 136768
rect 1258 134496 558742 135200
rect 1258 132928 558742 133632
rect 1258 131360 558742 132064
rect 1258 129792 558742 130496
rect 1258 128224 558742 128928
rect 1258 126656 558742 127360
rect 1258 125088 558742 125792
rect 1258 123520 558742 124224
rect 1258 121952 558742 122656
rect 1258 120384 558742 121088
rect 1258 118816 558742 119520
rect 1258 117248 558742 117952
rect 1258 115680 558742 116384
rect 1258 114112 558742 114816
rect 1258 112544 558742 113248
rect 1258 110976 558742 111680
rect 1258 109408 558742 110112
rect 1258 107840 558742 108544
rect 1258 106272 558742 106976
rect 1258 104704 558742 105408
rect 1258 103136 558742 103840
rect 1258 101568 558742 102272
rect 1258 100000 558742 100704
rect 1258 98432 558742 99136
rect 1258 96864 558742 97568
rect 1258 95296 558742 96000
rect 1258 93728 558742 94432
rect 1258 92160 558742 92864
rect 1258 90592 558742 91296
rect 1258 89024 558742 89728
rect 1258 87456 558742 88160
rect 1258 85888 558742 86592
rect 1258 84320 558742 85024
rect 1258 82752 558742 83456
rect 1258 81184 558742 81888
rect 1258 79616 558742 80320
rect 1258 78048 558742 78752
rect 1258 76480 558742 77184
rect 1258 74912 558742 75616
rect 1258 73344 558742 74048
rect 1258 71776 558742 72480
rect 1258 70208 558742 70912
rect 1258 68640 558742 69344
rect 1258 67072 558742 67776
rect 1258 65504 558742 66208
rect 1258 63936 558742 64640
rect 1258 62368 558742 63072
rect 1258 60800 558742 61504
rect 1258 59232 558742 59936
rect 1258 57664 558742 58368
rect 1258 56096 558742 56800
rect 1258 54528 558742 55232
rect 1258 52960 558742 53664
rect 1258 51392 558742 52096
rect 1258 49824 558742 50528
rect 1258 48256 558742 48960
rect 1258 46688 558742 47392
rect 1258 45120 558742 45824
rect 1258 43552 558742 44256
rect 1258 41984 558742 42688
rect 1258 40416 558742 41120
rect 1258 38848 558742 39552
rect 1258 37280 558742 37984
rect 1258 35712 558742 36416
rect 1258 34144 558742 34848
rect 1258 32576 558742 33280
rect 1258 31008 558742 31712
rect 1258 29440 558742 30144
rect 1258 27872 558742 28576
rect 1258 26304 558742 27008
rect 1258 24736 558742 25440
rect 1258 23168 558742 23872
rect 1258 21600 558742 22304
rect 1258 20032 558742 20736
rect 1258 18464 558742 19168
rect 1258 16896 558742 17600
rect 1258 15328 558742 16032
rect 1258 13760 558742 14464
rect 1258 12192 558742 12896
rect 1258 10624 558742 11328
rect 1258 9056 558742 9760
rect 1258 7488 558742 8192
rect 1258 5920 558742 6624
rect 1258 4352 558742 5056
rect 1258 3050 558742 3488
<< obsm1 >>
rect 1344 3076 558656 236828
<< metal2 >>
rect 263424 239200 263536 240000
rect 266784 239200 266896 240000
rect 290304 239200 290416 240000
rect 292320 239200 292432 240000
rect 300384 239200 300496 240000
rect 268800 0 268912 800
rect 269472 0 269584 800
rect 270144 0 270256 800
rect 270816 0 270928 800
rect 271488 0 271600 800
rect 272160 0 272272 800
rect 272832 0 272944 800
rect 274176 0 274288 800
rect 276864 0 276976 800
rect 281568 0 281680 800
rect 286272 0 286384 800
rect 287616 0 287728 800
rect 294336 0 294448 800
rect 309120 0 309232 800
rect 336000 0 336112 800
<< obsm2 >>
rect 4476 239140 263364 239200
rect 263596 239140 266724 239200
rect 266956 239140 290244 239200
rect 290476 239140 292260 239200
rect 292492 239140 300324 239200
rect 300556 239140 557700 239200
rect 4476 860 557700 239140
rect 4476 700 268740 860
rect 268972 700 269412 860
rect 269644 700 270084 860
rect 270316 700 270756 860
rect 270988 700 271428 860
rect 271660 700 272100 860
rect 272332 700 272772 860
rect 273004 700 274116 860
rect 274348 700 276804 860
rect 277036 700 281508 860
rect 281740 700 286212 860
rect 286444 700 287556 860
rect 287788 700 294276 860
rect 294508 700 309060 860
rect 309292 700 335940 860
rect 336172 700 557700 860
<< obsm3 >>
rect 4466 3108 557710 236796
<< metal4 >>
rect 4448 3076 4768 236828
rect 19808 3076 20128 236828
rect 35168 3076 35488 236828
rect 50528 3076 50848 236828
rect 65888 3076 66208 236828
rect 81248 3076 81568 236828
rect 96608 3076 96928 236828
rect 111968 3076 112288 236828
rect 127328 3076 127648 236828
rect 142688 3076 143008 236828
rect 158048 3076 158368 236828
rect 173408 3076 173728 236828
rect 188768 3076 189088 236828
rect 204128 3076 204448 236828
rect 219488 3076 219808 236828
rect 234848 3076 235168 236828
rect 250208 3076 250528 236828
rect 265568 3076 265888 236828
rect 280928 3076 281248 236828
rect 296288 3076 296608 236828
rect 311648 3076 311968 236828
rect 327008 3076 327328 236828
rect 342368 3076 342688 236828
rect 357728 3076 358048 236828
rect 373088 3076 373408 236828
rect 388448 3076 388768 236828
rect 403808 3076 404128 236828
rect 419168 3076 419488 236828
rect 434528 3076 434848 236828
rect 449888 3076 450208 236828
rect 465248 3076 465568 236828
rect 480608 3076 480928 236828
rect 495968 3076 496288 236828
rect 511328 3076 511648 236828
rect 526688 3076 527008 236828
rect 542048 3076 542368 236828
rect 557408 3076 557728 236828
<< obsm4 >>
rect 282156 113922 296228 119150
rect 296668 113922 298228 119150
<< labels >>
rlabel metal2 s 272832 0 272944 800 6 clk
port 1 nsew signal input
rlabel metal2 s 274176 0 274288 800 6 io_frequency[0]
port 2 nsew signal input
rlabel metal2 s 272160 0 272272 800 6 io_frequency[1]
port 3 nsew signal input
rlabel metal2 s 271488 0 271600 800 6 io_frequency[2]
port 4 nsew signal input
rlabel metal2 s 270144 0 270256 800 6 io_frequency[3]
port 5 nsew signal input
rlabel metal2 s 269472 0 269584 800 6 io_frequency[4]
port 6 nsew signal input
rlabel metal2 s 266784 239200 266896 240000 6 io_frequency[5]
port 7 nsew signal input
rlabel metal2 s 268800 0 268912 800 6 io_frequency[6]
port 8 nsew signal input
rlabel metal2 s 270816 0 270928 800 6 io_frequency[7]
port 9 nsew signal input
rlabel metal2 s 309120 0 309232 800 6 io_oeb_high[0]
port 10 nsew signal output
rlabel metal2 s 263424 239200 263536 240000 6 io_oeb_high[1]
port 11 nsew signal output
rlabel metal2 s 290304 239200 290416 240000 6 io_oeb_high[2]
port 12 nsew signal output
rlabel metal2 s 287616 0 287728 800 6 io_oeb_high[3]
port 13 nsew signal output
rlabel metal2 s 292320 239200 292432 240000 6 io_oeb_high[4]
port 14 nsew signal output
rlabel metal2 s 286272 0 286384 800 6 io_oeb_high[5]
port 15 nsew signal output
rlabel metal2 s 276864 0 276976 800 6 io_oeb_high[6]
port 16 nsew signal output
rlabel metal2 s 336000 0 336112 800 6 io_oeb_high[7]
port 17 nsew signal output
rlabel metal2 s 300384 239200 300496 240000 6 io_oeb_low
port 18 nsew signal output
rlabel metal2 s 294336 0 294448 800 6 io_pwm_1
port 19 nsew signal output
rlabel metal2 s 281568 0 281680 800 6 reset
port 20 nsew signal input
rlabel metal4 s 4448 3076 4768 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 526688 3076 527008 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 557408 3076 557728 236828 6 vdd
port 21 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 236828 6 vss
port 22 nsew ground bidirectional
rlabel metal4 s 542048 3076 542368 236828 6 vss
port 22 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 560000 240000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10998704
string GDS_FILE /home/moss/eda_tools_gf180_audiopwm/caravel_user_project/openlane/PWMaudio/runs/23_12_11_18_23/results/signoff/PWMaudio.magic.gds
string GDS_START 281950
<< end >>

