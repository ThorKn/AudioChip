VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO PWMaudio
  CLASS BLOCK ;
  FOREIGN PWMaudio ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 0.000 1388.240 4.000 ;
    END
  END clk
  PIN io_adsr_choice[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1323.840 1196.000 1324.400 1200.000 ;
    END
  END io_adsr_choice[0]
  PIN io_adsr_choice[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1327.200 1196.000 1327.760 1200.000 ;
    END
  END io_adsr_choice[1]
  PIN io_adsr_choice[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.480 1196.000 1321.040 1200.000 ;
    END
  END io_adsr_choice[2]
  PIN io_adsr_switch
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1428.000 0.000 1428.560 4.000 ;
    END
  END io_adsr_switch
  PIN io_frequency[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1377.600 0.000 1378.160 4.000 ;
    END
  END io_frequency[0]
  PIN io_frequency[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 0.000 1368.080 4.000 ;
    END
  END io_frequency[10]
  PIN io_frequency[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 0.000 1374.800 4.000 ;
    END
  END io_frequency[11]
  PIN io_frequency[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1370.880 0.000 1371.440 4.000 ;
    END
  END io_frequency[1]
  PIN io_frequency[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.960 0.000 1381.520 4.000 ;
    END
  END io_frequency[2]
  PIN io_frequency[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1364.160 0.000 1364.720 4.000 ;
    END
  END io_frequency[3]
  PIN io_frequency[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1360.800 0.000 1361.360 4.000 ;
    END
  END io_frequency[4]
  PIN io_frequency[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1350.720 0.000 1351.280 4.000 ;
    END
  END io_frequency[5]
  PIN io_frequency[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1357.440 0.000 1358.000 4.000 ;
    END
  END io_frequency[6]
  PIN io_frequency[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1344.000 0.000 1344.560 4.000 ;
    END
  END io_frequency[7]
  PIN io_frequency[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 0.000 1347.920 4.000 ;
    END
  END io_frequency[8]
  PIN io_frequency[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 0.000 1354.640 4.000 ;
    END
  END io_frequency[9]
  PIN io_loop
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1481.760 0.000 1482.320 4.000 ;
    END
  END io_loop
  PIN io_note_length[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 1196.000 1300.880 1200.000 ;
    END
  END io_note_length[0]
  PIN io_note_length[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 1196.000 1347.920 1200.000 ;
    END
  END io_note_length[1]
  PIN io_note_length[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1360.800 1196.000 1361.360 1200.000 ;
    END
  END io_note_length[2]
  PIN io_oeb_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1706.880 0.000 1707.440 4.000 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1438.080 0.000 1438.640 4.000 ;
    END
  END io_oeb_high[10]
  PIN io_oeb_high[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1612.800 0.000 1613.360 4.000 ;
    END
  END io_oeb_high[11]
  PIN io_oeb_high[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1535.520 0.000 1536.080 4.000 ;
    END
  END io_oeb_high[12]
  PIN io_oeb_high[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1552.320 1196.000 1552.880 1200.000 ;
    END
  END io_oeb_high[13]
  PIN io_oeb_high[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 0.000 1657.040 4.000 ;
    END
  END io_oeb_high[14]
  PIN io_oeb_high[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1643.040 1196.000 1643.600 1200.000 ;
    END
  END io_oeb_high[15]
  PIN io_oeb_high[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1656.480 1196.000 1657.040 1200.000 ;
    END
  END io_oeb_high[16]
  PIN io_oeb_high[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1088.640 0.000 1089.200 4.000 ;
    END
  END io_oeb_high[17]
  PIN io_oeb_high[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1676.640 0.000 1677.200 4.000 ;
    END
  END io_oeb_high[18]
  PIN io_oeb_high[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1464.960 1196.000 1465.520 1200.000 ;
    END
  END io_oeb_high[19]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1646.400 1196.000 1646.960 1200.000 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1438.080 1196.000 1438.640 1200.000 ;
    END
  END io_oeb_high[20]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1478.400 0.000 1478.960 4.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1404.480 0.000 1405.040 4.000 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1471.680 1196.000 1472.240 1200.000 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1317.120 0.000 1317.680 4.000 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1384.320 0.000 1384.880 4.000 ;
    END
  END io_oeb_high[6]
  PIN io_oeb_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1501.920 1196.000 1502.480 1200.000 ;
    END
  END io_oeb_high[7]
  PIN io_oeb_high[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1431.360 0.000 1431.920 4.000 ;
    END
  END io_oeb_high[8]
  PIN io_oeb_high[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 0.000 1556.240 4.000 ;
    END
  END io_oeb_high[9]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 1196.000 1354.640 1200.000 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1350.720 1196.000 1351.280 1200.000 ;
    END
  END io_oeb_low[1]
  PIN io_pwm_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.720 0.000 1435.280 4.000 ;
    END
  END io_pwm_1
  PIN io_pwm_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1475.040 0.000 1475.600 4.000 ;
    END
  END io_pwm_2
  PIN io_trigger
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1485.120 0.000 1485.680 4.000 ;
    END
  END io_trigger
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1401.120 0.000 1401.680 4.000 ;
    END
  END reset
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1184.140 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1184.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1184.140 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 1182.080 2793.710 1184.270 ;
      LAYER Nwell ;
        RECT 6.290 1177.760 2793.710 1182.080 ;
      LAYER Pwell ;
        RECT 6.290 1174.240 2793.710 1177.760 ;
      LAYER Nwell ;
        RECT 6.290 1169.920 2793.710 1174.240 ;
      LAYER Pwell ;
        RECT 6.290 1166.400 2793.710 1169.920 ;
      LAYER Nwell ;
        RECT 6.290 1162.080 2793.710 1166.400 ;
      LAYER Pwell ;
        RECT 6.290 1158.560 2793.710 1162.080 ;
      LAYER Nwell ;
        RECT 6.290 1154.240 2793.710 1158.560 ;
      LAYER Pwell ;
        RECT 6.290 1150.720 2793.710 1154.240 ;
      LAYER Nwell ;
        RECT 6.290 1146.400 2793.710 1150.720 ;
      LAYER Pwell ;
        RECT 6.290 1142.880 2793.710 1146.400 ;
      LAYER Nwell ;
        RECT 6.290 1138.560 2793.710 1142.880 ;
      LAYER Pwell ;
        RECT 6.290 1135.040 2793.710 1138.560 ;
      LAYER Nwell ;
        RECT 6.290 1130.720 2793.710 1135.040 ;
      LAYER Pwell ;
        RECT 6.290 1127.200 2793.710 1130.720 ;
      LAYER Nwell ;
        RECT 6.290 1122.880 2793.710 1127.200 ;
      LAYER Pwell ;
        RECT 6.290 1119.360 2793.710 1122.880 ;
      LAYER Nwell ;
        RECT 6.290 1115.040 2793.710 1119.360 ;
      LAYER Pwell ;
        RECT 6.290 1111.520 2793.710 1115.040 ;
      LAYER Nwell ;
        RECT 6.290 1107.200 2793.710 1111.520 ;
      LAYER Pwell ;
        RECT 6.290 1103.680 2793.710 1107.200 ;
      LAYER Nwell ;
        RECT 6.290 1099.360 2793.710 1103.680 ;
      LAYER Pwell ;
        RECT 6.290 1095.840 2793.710 1099.360 ;
      LAYER Nwell ;
        RECT 6.290 1091.520 2793.710 1095.840 ;
      LAYER Pwell ;
        RECT 6.290 1088.000 2793.710 1091.520 ;
      LAYER Nwell ;
        RECT 6.290 1083.680 2793.710 1088.000 ;
      LAYER Pwell ;
        RECT 6.290 1080.160 2793.710 1083.680 ;
      LAYER Nwell ;
        RECT 6.290 1075.840 2793.710 1080.160 ;
      LAYER Pwell ;
        RECT 6.290 1072.320 2793.710 1075.840 ;
      LAYER Nwell ;
        RECT 6.290 1068.000 2793.710 1072.320 ;
      LAYER Pwell ;
        RECT 6.290 1064.480 2793.710 1068.000 ;
      LAYER Nwell ;
        RECT 6.290 1060.160 2793.710 1064.480 ;
      LAYER Pwell ;
        RECT 6.290 1056.640 2793.710 1060.160 ;
      LAYER Nwell ;
        RECT 6.290 1052.320 2793.710 1056.640 ;
      LAYER Pwell ;
        RECT 6.290 1048.800 2793.710 1052.320 ;
      LAYER Nwell ;
        RECT 6.290 1044.480 2793.710 1048.800 ;
      LAYER Pwell ;
        RECT 6.290 1040.960 2793.710 1044.480 ;
      LAYER Nwell ;
        RECT 6.290 1036.640 2793.710 1040.960 ;
      LAYER Pwell ;
        RECT 6.290 1033.120 2793.710 1036.640 ;
      LAYER Nwell ;
        RECT 6.290 1028.800 2793.710 1033.120 ;
      LAYER Pwell ;
        RECT 6.290 1025.280 2793.710 1028.800 ;
      LAYER Nwell ;
        RECT 6.290 1020.960 2793.710 1025.280 ;
      LAYER Pwell ;
        RECT 6.290 1017.440 2793.710 1020.960 ;
      LAYER Nwell ;
        RECT 6.290 1013.120 2793.710 1017.440 ;
      LAYER Pwell ;
        RECT 6.290 1009.600 2793.710 1013.120 ;
      LAYER Nwell ;
        RECT 6.290 1005.280 2793.710 1009.600 ;
      LAYER Pwell ;
        RECT 6.290 1001.760 2793.710 1005.280 ;
      LAYER Nwell ;
        RECT 6.290 997.440 2793.710 1001.760 ;
      LAYER Pwell ;
        RECT 6.290 993.920 2793.710 997.440 ;
      LAYER Nwell ;
        RECT 6.290 989.600 2793.710 993.920 ;
      LAYER Pwell ;
        RECT 6.290 986.080 2793.710 989.600 ;
      LAYER Nwell ;
        RECT 6.290 981.760 2793.710 986.080 ;
      LAYER Pwell ;
        RECT 6.290 978.240 2793.710 981.760 ;
      LAYER Nwell ;
        RECT 6.290 973.920 2793.710 978.240 ;
      LAYER Pwell ;
        RECT 6.290 970.400 2793.710 973.920 ;
      LAYER Nwell ;
        RECT 6.290 966.080 2793.710 970.400 ;
      LAYER Pwell ;
        RECT 6.290 962.560 2793.710 966.080 ;
      LAYER Nwell ;
        RECT 6.290 958.240 2793.710 962.560 ;
      LAYER Pwell ;
        RECT 6.290 954.720 2793.710 958.240 ;
      LAYER Nwell ;
        RECT 6.290 950.400 2793.710 954.720 ;
      LAYER Pwell ;
        RECT 6.290 946.880 2793.710 950.400 ;
      LAYER Nwell ;
        RECT 6.290 942.560 2793.710 946.880 ;
      LAYER Pwell ;
        RECT 6.290 939.040 2793.710 942.560 ;
      LAYER Nwell ;
        RECT 6.290 934.720 2793.710 939.040 ;
      LAYER Pwell ;
        RECT 6.290 931.200 2793.710 934.720 ;
      LAYER Nwell ;
        RECT 6.290 926.880 2793.710 931.200 ;
      LAYER Pwell ;
        RECT 6.290 923.360 2793.710 926.880 ;
      LAYER Nwell ;
        RECT 6.290 919.040 2793.710 923.360 ;
      LAYER Pwell ;
        RECT 6.290 915.520 2793.710 919.040 ;
      LAYER Nwell ;
        RECT 6.290 911.200 2793.710 915.520 ;
      LAYER Pwell ;
        RECT 6.290 907.680 2793.710 911.200 ;
      LAYER Nwell ;
        RECT 6.290 903.360 2793.710 907.680 ;
      LAYER Pwell ;
        RECT 6.290 899.840 2793.710 903.360 ;
      LAYER Nwell ;
        RECT 6.290 895.520 2793.710 899.840 ;
      LAYER Pwell ;
        RECT 6.290 892.000 2793.710 895.520 ;
      LAYER Nwell ;
        RECT 6.290 887.680 2793.710 892.000 ;
      LAYER Pwell ;
        RECT 6.290 884.160 2793.710 887.680 ;
      LAYER Nwell ;
        RECT 6.290 879.840 2793.710 884.160 ;
      LAYER Pwell ;
        RECT 6.290 876.320 2793.710 879.840 ;
      LAYER Nwell ;
        RECT 6.290 872.000 2793.710 876.320 ;
      LAYER Pwell ;
        RECT 6.290 868.480 2793.710 872.000 ;
      LAYER Nwell ;
        RECT 6.290 864.160 2793.710 868.480 ;
      LAYER Pwell ;
        RECT 6.290 860.640 2793.710 864.160 ;
      LAYER Nwell ;
        RECT 6.290 856.320 2793.710 860.640 ;
      LAYER Pwell ;
        RECT 6.290 852.800 2793.710 856.320 ;
      LAYER Nwell ;
        RECT 6.290 848.480 2793.710 852.800 ;
      LAYER Pwell ;
        RECT 6.290 844.960 2793.710 848.480 ;
      LAYER Nwell ;
        RECT 6.290 840.640 2793.710 844.960 ;
      LAYER Pwell ;
        RECT 6.290 837.120 2793.710 840.640 ;
      LAYER Nwell ;
        RECT 6.290 832.800 2793.710 837.120 ;
      LAYER Pwell ;
        RECT 6.290 829.280 2793.710 832.800 ;
      LAYER Nwell ;
        RECT 6.290 824.960 2793.710 829.280 ;
      LAYER Pwell ;
        RECT 6.290 821.440 2793.710 824.960 ;
      LAYER Nwell ;
        RECT 6.290 817.120 2793.710 821.440 ;
      LAYER Pwell ;
        RECT 6.290 813.600 2793.710 817.120 ;
      LAYER Nwell ;
        RECT 6.290 809.280 2793.710 813.600 ;
      LAYER Pwell ;
        RECT 6.290 805.760 2793.710 809.280 ;
      LAYER Nwell ;
        RECT 6.290 801.440 2793.710 805.760 ;
      LAYER Pwell ;
        RECT 6.290 797.920 2793.710 801.440 ;
      LAYER Nwell ;
        RECT 6.290 793.600 2793.710 797.920 ;
      LAYER Pwell ;
        RECT 6.290 790.080 2793.710 793.600 ;
      LAYER Nwell ;
        RECT 6.290 785.760 2793.710 790.080 ;
      LAYER Pwell ;
        RECT 6.290 782.240 2793.710 785.760 ;
      LAYER Nwell ;
        RECT 6.290 777.920 2793.710 782.240 ;
      LAYER Pwell ;
        RECT 6.290 774.400 2793.710 777.920 ;
      LAYER Nwell ;
        RECT 6.290 770.080 2793.710 774.400 ;
      LAYER Pwell ;
        RECT 6.290 766.560 2793.710 770.080 ;
      LAYER Nwell ;
        RECT 6.290 762.240 2793.710 766.560 ;
      LAYER Pwell ;
        RECT 6.290 758.720 2793.710 762.240 ;
      LAYER Nwell ;
        RECT 6.290 754.400 2793.710 758.720 ;
      LAYER Pwell ;
        RECT 6.290 750.880 2793.710 754.400 ;
      LAYER Nwell ;
        RECT 6.290 746.560 2793.710 750.880 ;
      LAYER Pwell ;
        RECT 6.290 743.040 2793.710 746.560 ;
      LAYER Nwell ;
        RECT 6.290 738.845 2793.710 743.040 ;
        RECT 6.290 738.720 1393.430 738.845 ;
      LAYER Pwell ;
        RECT 6.290 735.200 2793.710 738.720 ;
      LAYER Nwell ;
        RECT 6.290 735.075 1350.625 735.200 ;
        RECT 6.290 731.005 2793.710 735.075 ;
        RECT 6.290 730.880 1324.305 731.005 ;
      LAYER Pwell ;
        RECT 6.290 727.360 2793.710 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 1363.750 727.360 ;
        RECT 6.290 723.040 2793.710 727.235 ;
      LAYER Pwell ;
        RECT 6.290 719.520 2793.710 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 1292.350 719.520 ;
        RECT 6.290 715.325 2793.710 719.395 ;
        RECT 6.290 715.200 1283.435 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 2793.710 715.200 ;
      LAYER Nwell ;
        RECT 6.290 707.360 2793.710 711.680 ;
      LAYER Pwell ;
        RECT 6.290 703.840 2793.710 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 1412.970 703.840 ;
        RECT 6.290 699.645 2793.710 703.715 ;
        RECT 6.290 699.520 1314.785 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 2793.710 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 1269.950 696.000 ;
        RECT 6.290 691.805 2793.710 695.875 ;
        RECT 6.290 691.680 1367.540 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 2793.710 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 1273.030 688.160 ;
        RECT 6.290 683.965 2793.710 688.035 ;
        RECT 6.290 683.840 1273.345 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 2793.710 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 1371.030 680.320 ;
        RECT 6.290 676.125 2793.710 680.195 ;
        RECT 6.290 676.000 1282.975 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 2793.710 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 1303.035 672.480 ;
        RECT 6.290 668.285 2793.710 672.355 ;
        RECT 6.290 668.160 1463.145 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 2793.710 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 1275.830 664.640 ;
        RECT 6.290 660.455 2793.710 664.515 ;
        RECT 6.290 660.445 1491.920 660.455 ;
        RECT 6.290 660.320 1304.390 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 2793.710 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 1291.510 656.800 ;
        RECT 6.290 652.615 2793.710 656.675 ;
        RECT 6.290 652.605 1491.920 652.615 ;
        RECT 6.290 652.480 1417.925 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 2793.710 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 1385.345 648.960 ;
        RECT 6.290 644.765 2793.710 648.835 ;
        RECT 6.290 644.640 1299.350 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 2793.710 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 1297.110 641.120 ;
        RECT 6.290 636.935 2793.710 640.995 ;
        RECT 6.290 636.925 1498.080 636.935 ;
        RECT 6.290 636.800 1369.115 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 2793.710 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 1317.045 633.280 ;
        RECT 6.290 629.095 2793.710 633.155 ;
        RECT 6.290 628.960 1495.840 629.095 ;
      LAYER Pwell ;
        RECT 6.290 625.440 2793.710 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 1421.235 625.440 ;
        RECT 6.290 621.245 2793.710 625.315 ;
        RECT 6.290 621.120 1423.555 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 2793.710 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 1370.185 617.600 ;
        RECT 6.290 613.415 2793.710 617.475 ;
        RECT 6.290 613.405 1496.960 613.415 ;
        RECT 6.290 613.280 1378.870 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 2793.710 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.625 1323.360 609.760 ;
        RECT 6.290 605.575 2793.710 609.625 ;
        RECT 6.290 605.440 1410.160 605.575 ;
      LAYER Pwell ;
        RECT 6.290 601.920 2793.710 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.785 1320.000 601.920 ;
        RECT 6.290 597.600 2793.710 601.785 ;
      LAYER Pwell ;
        RECT 6.290 594.080 2793.710 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.945 1322.240 594.080 ;
        RECT 6.290 589.895 2793.710 593.945 ;
        RECT 6.290 589.760 1386.640 589.895 ;
      LAYER Pwell ;
        RECT 6.290 586.240 2793.710 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.105 1428.640 586.240 ;
        RECT 6.290 582.055 2793.710 586.105 ;
        RECT 6.290 581.920 1342.400 582.055 ;
      LAYER Pwell ;
        RECT 6.290 578.400 2793.710 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.265 1358.080 578.400 ;
        RECT 6.290 574.215 2793.710 578.265 ;
        RECT 6.290 574.080 1419.120 574.215 ;
      LAYER Pwell ;
        RECT 6.290 570.560 2793.710 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.425 1360.880 570.560 ;
        RECT 6.290 566.365 2793.710 570.425 ;
        RECT 6.290 566.240 1483.445 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 2793.710 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.585 1369.280 562.720 ;
        RECT 6.290 558.535 2793.710 562.585 ;
        RECT 6.290 558.400 1497.520 558.535 ;
      LAYER Pwell ;
        RECT 6.290 554.880 2793.710 558.400 ;
      LAYER Nwell ;
        RECT 6.290 550.695 2793.710 554.880 ;
        RECT 6.290 550.560 1414.080 550.695 ;
      LAYER Pwell ;
        RECT 6.290 547.040 2793.710 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.905 1367.040 547.040 ;
        RECT 6.290 542.855 2793.710 546.905 ;
        RECT 6.290 542.720 1369.840 542.855 ;
      LAYER Pwell ;
        RECT 6.290 539.200 2793.710 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.065 1397.280 539.200 ;
        RECT 6.290 535.015 2793.710 539.065 ;
        RECT 6.290 534.880 1419.120 535.015 ;
      LAYER Pwell ;
        RECT 6.290 531.360 2793.710 534.880 ;
      LAYER Nwell ;
        RECT 6.290 527.175 2793.710 531.360 ;
        RECT 6.290 527.040 1383.280 527.175 ;
      LAYER Pwell ;
        RECT 6.290 523.520 2793.710 527.040 ;
      LAYER Nwell ;
        RECT 6.290 519.335 2793.710 523.520 ;
        RECT 6.290 519.325 1506.480 519.335 ;
        RECT 6.290 519.200 1411.630 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 2793.710 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.545 1355.280 515.680 ;
        RECT 6.290 511.495 2793.710 515.545 ;
        RECT 6.290 511.360 1349.120 511.495 ;
      LAYER Pwell ;
        RECT 6.290 507.840 2793.710 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.705 1401.760 507.840 ;
        RECT 6.290 503.655 2793.710 507.705 ;
        RECT 6.290 503.520 1327.565 503.655 ;
      LAYER Pwell ;
        RECT 6.290 500.000 2793.710 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 1425.070 500.000 ;
        RECT 6.290 499.865 1479.040 499.875 ;
        RECT 6.290 495.815 2793.710 499.865 ;
        RECT 6.290 495.805 1418.560 495.815 ;
        RECT 6.290 495.680 1367.390 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 2793.710 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.025 1447.680 492.160 ;
        RECT 6.290 487.975 2793.710 492.025 ;
        RECT 6.290 487.840 1416.880 487.975 ;
      LAYER Pwell ;
        RECT 6.290 484.320 2793.710 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.185 1323.360 484.320 ;
        RECT 6.290 480.135 2793.710 484.185 ;
        RECT 6.290 480.000 1382.720 480.135 ;
      LAYER Pwell ;
        RECT 6.290 476.480 2793.710 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.345 1323.920 476.480 ;
        RECT 6.290 472.295 2793.710 476.345 ;
        RECT 6.290 472.160 1418.000 472.295 ;
      LAYER Pwell ;
        RECT 6.290 468.640 2793.710 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.505 1330.080 468.640 ;
        RECT 6.290 464.455 2793.710 468.505 ;
        RECT 6.290 464.320 1487.440 464.455 ;
      LAYER Pwell ;
        RECT 6.290 460.800 2793.710 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.665 1350.240 460.800 ;
        RECT 6.290 456.480 2793.710 460.665 ;
      LAYER Pwell ;
        RECT 6.290 452.960 2793.710 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.825 1471.760 452.960 ;
        RECT 6.290 448.775 2793.710 452.825 ;
        RECT 6.290 448.640 1409.040 448.775 ;
      LAYER Pwell ;
        RECT 6.290 445.120 2793.710 448.640 ;
      LAYER Nwell ;
        RECT 6.290 440.800 2793.710 445.120 ;
      LAYER Pwell ;
        RECT 6.290 437.280 2793.710 440.800 ;
      LAYER Nwell ;
        RECT 6.290 432.960 2793.710 437.280 ;
      LAYER Pwell ;
        RECT 6.290 429.440 2793.710 432.960 ;
      LAYER Nwell ;
        RECT 6.290 425.120 2793.710 429.440 ;
      LAYER Pwell ;
        RECT 6.290 421.600 2793.710 425.120 ;
      LAYER Nwell ;
        RECT 6.290 417.280 2793.710 421.600 ;
      LAYER Pwell ;
        RECT 6.290 413.760 2793.710 417.280 ;
      LAYER Nwell ;
        RECT 6.290 409.440 2793.710 413.760 ;
      LAYER Pwell ;
        RECT 6.290 405.920 2793.710 409.440 ;
      LAYER Nwell ;
        RECT 6.290 401.600 2793.710 405.920 ;
      LAYER Pwell ;
        RECT 6.290 398.080 2793.710 401.600 ;
      LAYER Nwell ;
        RECT 6.290 393.760 2793.710 398.080 ;
      LAYER Pwell ;
        RECT 6.290 390.240 2793.710 393.760 ;
      LAYER Nwell ;
        RECT 6.290 385.920 2793.710 390.240 ;
      LAYER Pwell ;
        RECT 6.290 382.400 2793.710 385.920 ;
      LAYER Nwell ;
        RECT 6.290 378.080 2793.710 382.400 ;
      LAYER Pwell ;
        RECT 6.290 374.560 2793.710 378.080 ;
      LAYER Nwell ;
        RECT 6.290 370.240 2793.710 374.560 ;
      LAYER Pwell ;
        RECT 6.290 366.720 2793.710 370.240 ;
      LAYER Nwell ;
        RECT 6.290 362.400 2793.710 366.720 ;
      LAYER Pwell ;
        RECT 6.290 358.880 2793.710 362.400 ;
      LAYER Nwell ;
        RECT 6.290 354.560 2793.710 358.880 ;
      LAYER Pwell ;
        RECT 6.290 351.040 2793.710 354.560 ;
      LAYER Nwell ;
        RECT 6.290 346.720 2793.710 351.040 ;
      LAYER Pwell ;
        RECT 6.290 343.200 2793.710 346.720 ;
      LAYER Nwell ;
        RECT 6.290 338.880 2793.710 343.200 ;
      LAYER Pwell ;
        RECT 6.290 335.360 2793.710 338.880 ;
      LAYER Nwell ;
        RECT 6.290 331.040 2793.710 335.360 ;
      LAYER Pwell ;
        RECT 6.290 327.520 2793.710 331.040 ;
      LAYER Nwell ;
        RECT 6.290 323.200 2793.710 327.520 ;
      LAYER Pwell ;
        RECT 6.290 319.680 2793.710 323.200 ;
      LAYER Nwell ;
        RECT 6.290 315.360 2793.710 319.680 ;
      LAYER Pwell ;
        RECT 6.290 311.840 2793.710 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.520 2793.710 311.840 ;
      LAYER Pwell ;
        RECT 6.290 304.000 2793.710 307.520 ;
      LAYER Nwell ;
        RECT 6.290 299.680 2793.710 304.000 ;
      LAYER Pwell ;
        RECT 6.290 296.160 2793.710 299.680 ;
      LAYER Nwell ;
        RECT 6.290 291.840 2793.710 296.160 ;
      LAYER Pwell ;
        RECT 6.290 288.320 2793.710 291.840 ;
      LAYER Nwell ;
        RECT 6.290 284.000 2793.710 288.320 ;
      LAYER Pwell ;
        RECT 6.290 280.480 2793.710 284.000 ;
      LAYER Nwell ;
        RECT 6.290 276.160 2793.710 280.480 ;
      LAYER Pwell ;
        RECT 6.290 272.640 2793.710 276.160 ;
      LAYER Nwell ;
        RECT 6.290 268.320 2793.710 272.640 ;
      LAYER Pwell ;
        RECT 6.290 264.800 2793.710 268.320 ;
      LAYER Nwell ;
        RECT 6.290 260.480 2793.710 264.800 ;
      LAYER Pwell ;
        RECT 6.290 256.960 2793.710 260.480 ;
      LAYER Nwell ;
        RECT 6.290 252.640 2793.710 256.960 ;
      LAYER Pwell ;
        RECT 6.290 249.120 2793.710 252.640 ;
      LAYER Nwell ;
        RECT 6.290 244.800 2793.710 249.120 ;
      LAYER Pwell ;
        RECT 6.290 241.280 2793.710 244.800 ;
      LAYER Nwell ;
        RECT 6.290 236.960 2793.710 241.280 ;
      LAYER Pwell ;
        RECT 6.290 233.440 2793.710 236.960 ;
      LAYER Nwell ;
        RECT 6.290 229.120 2793.710 233.440 ;
      LAYER Pwell ;
        RECT 6.290 225.600 2793.710 229.120 ;
      LAYER Nwell ;
        RECT 6.290 221.280 2793.710 225.600 ;
      LAYER Pwell ;
        RECT 6.290 217.760 2793.710 221.280 ;
      LAYER Nwell ;
        RECT 6.290 213.440 2793.710 217.760 ;
      LAYER Pwell ;
        RECT 6.290 209.920 2793.710 213.440 ;
      LAYER Nwell ;
        RECT 6.290 205.600 2793.710 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 2793.710 205.600 ;
      LAYER Nwell ;
        RECT 6.290 197.760 2793.710 202.080 ;
      LAYER Pwell ;
        RECT 6.290 194.240 2793.710 197.760 ;
      LAYER Nwell ;
        RECT 6.290 189.920 2793.710 194.240 ;
      LAYER Pwell ;
        RECT 6.290 186.400 2793.710 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.080 2793.710 186.400 ;
      LAYER Pwell ;
        RECT 6.290 178.560 2793.710 182.080 ;
      LAYER Nwell ;
        RECT 6.290 174.240 2793.710 178.560 ;
      LAYER Pwell ;
        RECT 6.290 170.720 2793.710 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 2793.710 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 2793.710 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 2793.710 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 2793.710 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 2793.710 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 2793.710 150.720 ;
      LAYER Nwell ;
        RECT 6.290 142.880 2793.710 147.200 ;
      LAYER Pwell ;
        RECT 6.290 139.360 2793.710 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 2793.710 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 2793.710 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 2793.710 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 2793.710 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 2793.710 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 2793.710 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 2793.710 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 2793.710 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 2793.710 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 2793.710 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 2793.710 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 2793.710 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 2793.710 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 2793.710 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 2793.710 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 2793.710 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 2793.710 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 2793.710 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 2793.710 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 2793.710 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 2793.710 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 2793.710 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 2793.710 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 2793.710 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 2793.710 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 2793.710 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 2793.710 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 2793.710 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 2793.710 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 2793.710 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 2793.710 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 2793.710 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 14.710 2793.280 1184.140 ;
      LAYER Metal2 ;
        RECT 22.380 1195.700 1300.020 1196.000 ;
        RECT 1301.180 1195.700 1320.180 1196.000 ;
        RECT 1321.340 1195.700 1323.540 1196.000 ;
        RECT 1324.700 1195.700 1326.900 1196.000 ;
        RECT 1328.060 1195.700 1347.060 1196.000 ;
        RECT 1348.220 1195.700 1350.420 1196.000 ;
        RECT 1351.580 1195.700 1353.780 1196.000 ;
        RECT 1354.940 1195.700 1360.500 1196.000 ;
        RECT 1361.660 1195.700 1437.780 1196.000 ;
        RECT 1438.940 1195.700 1464.660 1196.000 ;
        RECT 1465.820 1195.700 1471.380 1196.000 ;
        RECT 1472.540 1195.700 1501.620 1196.000 ;
        RECT 1502.780 1195.700 1552.020 1196.000 ;
        RECT 1553.180 1195.700 1642.740 1196.000 ;
        RECT 1643.900 1195.700 1646.100 1196.000 ;
        RECT 1647.260 1195.700 1656.180 1196.000 ;
        RECT 1657.340 1195.700 2788.500 1196.000 ;
        RECT 22.380 4.300 2788.500 1195.700 ;
        RECT 22.380 3.500 1088.340 4.300 ;
        RECT 1089.500 3.500 1316.820 4.300 ;
        RECT 1317.980 3.500 1343.700 4.300 ;
        RECT 1344.860 3.500 1347.060 4.300 ;
        RECT 1348.220 3.500 1350.420 4.300 ;
        RECT 1351.580 3.500 1353.780 4.300 ;
        RECT 1354.940 3.500 1357.140 4.300 ;
        RECT 1358.300 3.500 1360.500 4.300 ;
        RECT 1361.660 3.500 1363.860 4.300 ;
        RECT 1365.020 3.500 1367.220 4.300 ;
        RECT 1368.380 3.500 1370.580 4.300 ;
        RECT 1371.740 3.500 1373.940 4.300 ;
        RECT 1375.100 3.500 1377.300 4.300 ;
        RECT 1378.460 3.500 1380.660 4.300 ;
        RECT 1381.820 3.500 1384.020 4.300 ;
        RECT 1385.180 3.500 1387.380 4.300 ;
        RECT 1388.540 3.500 1400.820 4.300 ;
        RECT 1401.980 3.500 1404.180 4.300 ;
        RECT 1405.340 3.500 1427.700 4.300 ;
        RECT 1428.860 3.500 1431.060 4.300 ;
        RECT 1432.220 3.500 1434.420 4.300 ;
        RECT 1435.580 3.500 1437.780 4.300 ;
        RECT 1438.940 3.500 1474.740 4.300 ;
        RECT 1475.900 3.500 1478.100 4.300 ;
        RECT 1479.260 3.500 1481.460 4.300 ;
        RECT 1482.620 3.500 1484.820 4.300 ;
        RECT 1485.980 3.500 1535.220 4.300 ;
        RECT 1536.380 3.500 1555.380 4.300 ;
        RECT 1556.540 3.500 1612.500 4.300 ;
        RECT 1613.660 3.500 1656.180 4.300 ;
        RECT 1657.340 3.500 1676.340 4.300 ;
        RECT 1677.500 3.500 1706.580 4.300 ;
        RECT 1707.740 3.500 2788.500 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 15.540 2788.550 1183.980 ;
      LAYER Metal4 ;
        RECT 1330.700 589.770 1404.340 718.390 ;
        RECT 1406.540 589.770 1481.140 718.390 ;
        RECT 1483.340 589.770 1486.660 718.390 ;
  END
END PWMaudio
END LIBRARY

